module tx_handshake_t.v();
   
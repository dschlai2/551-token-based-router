module tx_handshake_t();
   reg rc_has_data, 